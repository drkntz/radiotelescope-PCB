** Profile: "SCHEMATIC1-hbridge"  [ s:\projects\radiotelescope\radiotelescope-pcb\simulation\hbridge\hbridge-pspicefiles\schematic1\hbridge.sim ] 

** Creating circuit file "hbridge.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../hbridge-pspicefiles/hbridge.lib" 
* From [PSPICE NETLIST] section of C:\Users\zach\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 500u 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
